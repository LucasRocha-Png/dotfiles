context IEEE_BIT_CONTEXT is
  library IEEE;
  use IEEE.numeric_bit.all;
end context IEEE_BIT_CONTEXT;

context IEEE_STD_CONTEXT is
  library IEEE;
  use IEEE.std_logic_1164.all;
  use IEEE.Numeric_Std.all;
end context IEEE_STD_CONTEXT;