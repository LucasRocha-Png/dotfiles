-- Here you can try the package and/or entity-architecture snippets.
-- Just type 'pkgfull-' or 'entarch-'. While you start typing, a list of available snippets 
-- will pop up automatically. Choose the one you want and see what happens.

